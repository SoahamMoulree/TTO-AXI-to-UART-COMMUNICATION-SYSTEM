`define num_of_txns 8
`define baud_count 434
